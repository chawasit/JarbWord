module FinalBox();


endmodule
